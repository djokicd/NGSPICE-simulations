* Fast impulse diode, shows trr, ts

Vg 1 0 PULSE(0 1 2n 1p 1p 100n 200n 0)
R1 1 2 0.5k
D1 2 0 1N4148

.model 1N4148 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n Iave=200m Vpk=75)

.control
save all
tran 0.01n 1000n 0n
plot v(1) v(2)
plot -i(Vg)
