* Buffered current mirror ckt

.include bc337.ckt

I0 0 1 1m
Q1 1 2 0 bc337
Q2 3 2 0 bc337
Rshort1 3 2 0
Q3 4 1 3 bc337
Vout 4 0 2.5

* Output current into 4

.model generic npn

.control
save all @Q1[ib] @Q2[ib] @Q3[ib] @Q1[ic] @Q2[ic] @Q3[ic]
dc Vout 0.0 5.0 0.01
run
plot @Q1[ib] @Q2[ib] @Q3[ib]
plot @Q1[ic] @Q2[ic] @Q3[ic]

tf i(Vout) Vout
run
print transfer_function
